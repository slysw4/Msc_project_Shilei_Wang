module Rom(
	input wire clk,
	input wire [9:0] addr,
	
	output reg[2:0] weight1,
	output reg[2:0] weight2,
	output reg[2:0] weight3
);

reg [2:0] rom [287:0];

initial begin 

 rom [ 0  ]<= 3'd0;
 rom [ 1  ]<= 3'd0;
 rom [ 2  ]<= 3'd0;
 rom [ 3  ]<= 3'd0;
 rom [ 4  ]<= 3'd1;
 rom [ 5  ]<= 3'd0;
 rom [ 6  ]<= 3'd0;
 rom [ 7  ]<= 3'd0;
 rom [ 8  ]<= 3'd1;
 rom [ 9  ]<= 3'd2;
 rom [ 10  ]<= 3'd1;
 rom [ 11  ]<= 3'd0;
 rom [ 12  ]<= 3'd0;
 rom [ 13  ]<= 3'd0;
 rom [ 14  ]<= 3'd0;
 rom [ 15  ]<= 3'd1;
 rom [ 16  ]<= 3'd0;
 rom [ 17  ]<= 3'd0;
 rom [ 18  ]<= 3'd0;
 rom [ 19  ]<= 3'd0;
 rom [ 20  ]<= 3'd0;
 rom [ 21  ]<= 3'd0;
 rom [ 22  ]<= 3'd0;
 rom [ 23  ]<= 3'd0;
 rom [ 24  ]<= 3'd0;
 rom [ 25  ]<= 3'd0;
 rom [ 26  ]<= 3'd0;
 rom [ 27  ]<= 3'd0;
 rom [ 28  ]<= 3'd0;
 rom [ 29  ]<= 3'd0;
 rom [ 30  ]<= 3'd0;
 rom [ 31  ]<= 3'd0;
 rom [ 32  ]<= 3'd0;
 rom [ 33  ]<= 3'd0;
 rom [ 34  ]<= 3'd0;
 rom [ 35  ]<= 3'd0;
 rom [ 36  ]<= 3'd0;
 rom [ 37  ]<= 3'd0;
 rom [ 38  ]<= 3'd0;
 rom [ 39  ]<= 3'd0;
 rom [ 40  ]<= 3'd0;
 rom [ 41  ]<= 3'd0;
 rom [ 42  ]<= 3'd0;
 rom [ 43  ]<= 3'd0;
 rom [ 44  ]<= 3'd0;
 rom [ 45  ]<= 3'd0;
 rom [ 46  ]<= 3'd1;
 rom [ 47  ]<= 3'd1;
 rom [ 48  ]<= 3'd0;
 rom [ 49  ]<= 3'd1;
 rom [ 50  ]<= 3'd0;
 rom [ 51  ]<= 3'd0;
 rom [ 52  ]<= 3'd0;
 rom [ 53  ]<= 3'd0;
 rom [ 54  ]<= 3'd0;
 rom [ 55  ]<= 3'd0;
 rom [ 56  ]<= 3'd0;
 rom [ 57  ]<= 3'd0;
 rom [ 58  ]<= 3'd0;
 rom [ 59  ]<= 3'd0;
 rom [ 60  ]<= 3'd0;
 rom [ 61  ]<= 3'd0;
 rom [ 62  ]<= 3'd0;
 rom [ 63  ]<= 3'd0;
 rom [ 64  ]<= 3'd0;
 rom [ 65  ]<= 3'd0;
 rom [ 66  ]<= 3'd0;
 rom [ 67  ]<= 3'd0;
 rom [ 68  ]<= 3'd0;
 rom [ 69  ]<= 3'd0;
 rom [ 70  ]<= 3'd0;
 rom [ 71  ]<= 3'd0;
 rom [ 72  ]<= 3'd0;
 rom [ 73  ]<= 3'd0;
 rom [ 74  ]<= 3'd0;
 rom [ 75  ]<= 3'd0;
 rom [ 76  ]<= 3'd0;
 rom [ 77  ]<= 3'd0;
 rom [ 78  ]<= 3'd0;
 rom [ 79  ]<= 3'd0;
 rom [ 80  ]<= 3'd0;
 rom [ 81  ]<= 3'd0;
 rom [ 82  ]<= 3'd0;
 rom [ 83  ]<= 3'd0;
 rom [ 84  ]<= 3'd0;
 rom [ 85  ]<= 3'd0;
 rom [ 86  ]<= 3'd0;
 rom [ 87  ]<= 3'd0;
 rom [ 88  ]<= 3'd0;
 rom [ 89  ]<= 3'd0;
 rom [ 90  ]<= 3'd1;
 rom [ 91  ]<= 3'd0;
 rom [ 92  ]<= 3'd0;
 rom [ 93  ]<= 3'd0;
 rom [ 94  ]<= 3'd0;
 rom [ 95  ]<= 3'd0;
 rom [ 96  ]<= 3'd0;
 rom [ 97  ]<= 3'd0;
 rom [ 98  ]<= 3'd0;
 rom [ 99  ]<= 3'd0;
 rom [ 100  ]<= 3'd0;
 rom [ 101  ]<= 3'd0;
 rom [ 102  ]<= 3'd0;
 rom [ 103  ]<= 3'd0;
 rom [ 104  ]<= 3'd1;
 rom [ 105  ]<= 3'd1;
 rom [ 106  ]<= 3'd0;
 rom [ 107  ]<= 3'd0;
 rom [ 108  ]<= 3'd0;
 rom [ 109  ]<= 3'd0;
 rom [ 110  ]<= 3'd0;
 rom [ 111  ]<= 3'd0;
 rom [ 112  ]<= 3'd0;
 rom [ 113  ]<= 3'd0;
 rom [ 114  ]<= 3'd0;
 rom [ 115  ]<= 3'd0;
 rom [ 116  ]<= 3'd0;
 rom [ 117  ]<= 3'd0;
 rom [ 118  ]<= 3'd0;
 rom [ 119  ]<= 3'd0;
 rom [ 120  ]<= 3'd0;
 rom [ 121  ]<= 3'd0;
 rom [ 122  ]<= 3'd0;
 rom [ 123  ]<= 3'd0;
 rom [ 124  ]<= 3'd0;
 rom [ 125  ]<= 3'd0;
 rom [ 126  ]<= 3'd0;
 rom [ 127  ]<= 3'd0;
 rom [ 128  ]<= 3'd0;
 rom [ 129  ]<= 3'd0;
 rom [ 130  ]<= 3'd0;
 rom [ 131  ]<= 3'd0;
 rom [ 132  ]<= 3'd0;
 rom [ 133  ]<= 3'd0;
 rom [ 134  ]<= 3'd0;
 rom [ 135  ]<= 3'd0;
 rom [ 136  ]<= 3'd0;
 rom [ 137  ]<= 3'd0;
 rom [ 138  ]<= 3'd0;
 rom [ 139  ]<= 3'd0;
 rom [ 140  ]<= 3'd0;
 rom [ 141  ]<= 3'd0;
 rom [ 142  ]<= 3'd0;
 rom [ 143  ]<= 3'd0;
 rom [ 144  ]<= 3'd0;
 rom [ 145  ]<= 3'd0;
 rom [ 146  ]<= 3'd0;
 rom [ 147  ]<= 3'd0;
 rom [ 148  ]<= 3'd0;
 rom [ 149  ]<= 3'd0;
 rom [ 150  ]<= 3'd0;
 rom [ 151  ]<= 3'd0;
 rom [ 152  ]<= 3'd0;
 rom [ 153  ]<= 3'd0;
 rom [ 154  ]<= 3'd0;
 rom [ 155  ]<= 3'd0;
 rom [ 156  ]<= 3'd0;
 rom [ 157  ]<= 3'd0;
 rom [ 158  ]<= 3'd0;
 rom [ 159  ]<= 3'd0;
 rom [ 160  ]<= 3'd0;
 rom [ 161  ]<= 3'd0;
 rom [ 162  ]<= 3'd0;
 rom [ 163  ]<= 3'd0;
 rom [ 164  ]<= 3'd0;
 rom [ 165  ]<= 3'd0;
 rom [ 166  ]<= 3'd0;
 rom [ 167  ]<= 3'd0;
 rom [ 168  ]<= 3'd0;
 rom [ 169  ]<= 3'd0;
 rom [ 170  ]<= 3'd0;
 rom [ 171  ]<= 3'd0;
 rom [ 172  ]<= 3'd0;
 rom [ 173  ]<= 3'd0;
 rom [ 174  ]<= 3'd0;
 rom [ 175  ]<= 3'd0;
 rom [ 176  ]<= 3'd0;
 rom [ 177  ]<= 3'd0;
 rom [ 178  ]<= 3'd0;
 rom [ 179  ]<= 3'd0;
 rom [ 180  ]<= 3'd0;
 rom [ 181  ]<= 3'd0;
 rom [ 182  ]<= 3'd0;
 rom [ 183  ]<= 3'd0;
 rom [ 184  ]<= 3'd0;
 rom [ 185  ]<= 3'd0;
 rom [ 186  ]<= 3'd1;
 rom [ 187  ]<= 3'd0;
 rom [ 188  ]<= 3'd0;
 rom [ 189  ]<= 3'd0;
 rom [ 190  ]<= 3'd0;
 rom [ 191  ]<= 3'd0;
 rom [ 192  ]<= 3'd0;
 rom [ 193  ]<= 3'd0;
 rom [ 194  ]<= 3'd0;
 rom [ 195  ]<= 3'd0;
 rom [ 196  ]<= 3'd0;
 rom [ 197  ]<= 3'd0;
 rom [ 198  ]<= 3'd0;
 rom [ 199  ]<= 3'd0;
 rom [ 200  ]<= 3'd0;
 rom [ 201  ]<= 3'd0;
 rom [ 202  ]<= 3'd0;
 rom [ 203  ]<= 3'd0;
 rom [ 204  ]<= 3'd0;
 rom [ 205  ]<= 3'd0;
 rom [ 206  ]<= 3'd0;
 rom [ 207  ]<= 3'd0;
 rom [ 208  ]<= 3'd0;
 rom [ 209  ]<= 3'd0;
 rom [ 210  ]<= 3'd0;
 rom [ 211  ]<= 3'd0;
 rom [ 212  ]<= 3'd0;
 rom [ 213  ]<= 3'd0;
 rom [ 214  ]<= 3'd0;
 rom [ 215  ]<= 3'd0;
 rom [ 216  ]<= 3'd0;
 rom [ 217  ]<= 3'd0;
 rom [ 218  ]<= 3'd0;
 rom [ 219  ]<= 3'd0;
 rom [ 220  ]<= 3'd0;
 rom [ 221  ]<= 3'd0;
 rom [ 222  ]<= 3'd0;
 rom [ 223  ]<= 3'd0;
 rom [ 224  ]<= 3'd0;
 rom [ 225  ]<= 3'd0;
 rom [ 226  ]<= 3'd0;
 rom [ 227  ]<= 3'd0;
 rom [ 228  ]<= 3'd0;
 rom [ 229  ]<= 3'd0;
 rom [ 230  ]<= 3'd0;
 rom [ 231  ]<= 3'd0;
 rom [ 232  ]<= 3'd0;
 rom [ 233  ]<= 3'd0;
 rom [ 234  ]<= 3'd0;
 rom [ 235  ]<= 3'd0;
 rom [ 236  ]<= 3'd0;
 rom [ 237  ]<= 3'd0;
 rom [ 238  ]<= 3'd0;
 rom [ 239  ]<= 3'd0;
 rom [ 240  ]<= 3'd0;
 rom [ 241  ]<= 3'd0;
 rom [ 242  ]<= 3'd0;
 rom [ 243  ]<= 3'd0;
 rom [ 244  ]<= 3'd0;
 rom [ 245  ]<= 3'd0;
 rom [ 246  ]<= 3'd0;
 rom [ 247  ]<= 3'd0;
 rom [ 248  ]<= 3'd0;
 rom [ 249  ]<= 3'd0;
 rom [ 250  ]<= 3'd0;
 rom [ 251  ]<= 3'd0;
 rom [ 252  ]<= 3'd0;
 rom [ 253  ]<= 3'd0;
 rom [ 254  ]<= 3'd0;
 rom [ 255  ]<= 3'd0;
 rom [ 256  ]<= 3'd0;
 rom [ 257  ]<= 3'd0;
 rom [ 258  ]<= 3'd0;
 rom [ 259  ]<= 3'd0;
 rom [ 260  ]<= 3'd0;
 rom [ 261  ]<= 3'd0;
 rom [ 262  ]<= 3'd0;
 rom [ 263  ]<= 3'd0;
 rom [ 264  ]<= 3'd0;
 rom [ 265  ]<= 3'd0;
 rom [ 266  ]<= 3'd0;
 rom [ 267  ]<= 3'd0;
 rom [ 268  ]<= 3'd0;
 rom [ 269  ]<= 3'd0;
 rom [ 270  ]<= 3'd0;
 rom [ 271  ]<= 3'd0;
 rom [ 272  ]<= 3'd0;
 rom [ 273  ]<= 3'd0;
 rom [ 274  ]<= 3'd0;
 rom [ 275  ]<= 3'd0;
 rom [ 276  ]<= 3'd0;
 rom [ 277  ]<= 3'd0;
 rom [ 278  ]<= 3'd0;
 rom [ 279  ]<= 3'd0;
 rom [ 280  ]<= 3'd0;
 rom [ 281  ]<= 3'd0;
 rom [ 282  ]<= 3'd0;
 rom [ 283  ]<= 3'd0;
 rom [ 284  ]<= 3'd0;
 rom [ 285  ]<= 3'd0;
 rom [ 286  ]<= 3'd0;
 rom [ 287  ]<= 3'd0;

 
end


always@(posedge clk)
begin 
	weight1 <= rom[addr];
	weight2 <= rom[addr + 96];
	weight3 <= rom[addr + 192];
	end 
endmodule
